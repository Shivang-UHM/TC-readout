
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY GRAY_ENCODER IS
	GENERIC (
		NBITS : INTEGER := 8
	);
	PORT (
		GRAY_OUT : OUT STD_LOGIC_VECTOR(NBITS - 1 DOWNTO 0);
		BIN_IN : IN STD_LOGIC_VECTOR(NBITS - 1 DOWNTO 0)
	);
END GRAY_ENCODER;

ARCHITECTURE Behavioral OF GRAY_ENCODER IS

BEGIN

	GRAY_OUT(NBITS - 1) <= BIN_IN(NBITS - 1);

	GEN_XOR : FOR I IN 0 TO NBITS - 2 GENERATE
		GRAY_OUT(I) <= BIN_IN(I + 1) XOR BIN_IN(I);

	END GENERATE;

END Behavioral;